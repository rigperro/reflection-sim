0:(217,171):174
0:(307,247):215
2:(217,296):211
1:(835,404):113
0:(756,675):250
2:(772,180):265
1:(725,107):179
1:(815,382):252
3:(115,688):75
0:(114,524):196
0:(845,604):316
2:(683,479):128
2:(778,654):83
1:(422,198):253
2:(379,735):72
1:(898,636):161
3:(181,21):226
3:(152,55):298
0:(414,143):332
2:(196,144):321
1:(58,87):29
1:(354,50):314
1:(549,711):96
0:(148,109):105
0:(828,722):232
2:(770,561):265
3:(872,324):290
3:(302,459):55
3:(871,618):81
0:(715,28):279
2:(101,548):70
0:(537,365):207
0:(815,157):250
1:(60,760):63
1:(644,8):57
0:(407,475):306
1:(490,244):138
3:(604,785):354
1:(14,640):93
1:(582,182):234
1:(304,222):226
2:(3,228):168
0:(89,288):107
0:(168,720):327
1:(462,144):153
0:(887,364):234
0:(460,389):76
1:(136,395):21
#
